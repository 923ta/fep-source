DEMO CIRCUIT

.include 'LMC6482A.LIB'

.global vcc vee
vcc vcc 0 50
vee vee 0 -50

.ic v(7)=0v v(8)=0v v(9)=0v v(10)=0v v(11)=0v v(12)=0v v(13)=0v v(14)=0v v(15)=0v v(16)=0v v(17)=0v v(18)=0v v(19)=0v v(20)=0v v(21)=0v v(22)=0v

* εu,1 積分
x1 0 7 vcc vee 13 LMC6482A/NS
r1 1 7 100k
c1 7 13 100n

* εu,2 積分
x2 0 8 vcc vee 14 LMC6482A/NS
r2 2 8 100k
c2 8 14 100n

* φ1 積分
x3 0 9 vcc vee 15 LMC6482A/NS
r3 3 9 100k
c3 9 15 100n

* φ2 積分
x4 0 10 vcc vee 16 LMC6482A/NS
r4 4 10 100k
c4 10 16 100n

* εp,1 積分
x5 0 11 vcc vee 17 LMC6482A/NS
r5 5 11 100k
c5 11 17 100n

* εp,2 積分
x6 0 12 vcc vee 18 LMC6482A/NS
r6 6 12 100k
c6 12 18 100n

* φ1 反転
x7 0 19 vcc vee 21 LMC6482A/NS
r71 15 19 100k
r72 19 21 100k

* φ2 反転
x8 0 20 vcc vee 22 LMC6482A/NS
r81 16 20 100k
r82 20 22 100k

v1 23 0 1
v2 0 24 1
vu1 0 25 5
vu2 0 26 5

r11 13 1 100k ; Σu11
r12 14 1 100k ; Σu12
r13 15 1 101k ; θ11
r14 16 1 99k ; θ12
r15 25 1 100k
r16 13 2 100k ; Σu12
r17 14 2 100k ; Σu22
r18 15 2 99k ; θ21
r19 16 2 100k ; θ22
r20 26 2 100k
r21 17 3 100k
r22 24 3 100k ; θ11
r23 18 4 100k
r24 24 4 100k ; θ12
r25 21 5 100k
r26 17 5 100k ; Σp11
r27 18 5 100k ; Σp12
r28 23 5 25k ; vp1
r29 22 6 100k
r30 17 6 100k ; Σp12
r31 18 6 100k ; Σp22
r32 23 6 50k ; vp2

.control
tran 100u 10
plot v(13) v(14) v(17) v(18)
plot v(15) v(16)
.endc

.end