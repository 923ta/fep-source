DEMO CIRCUIT
* 関数g(φ)がφ^2 抵抗の単位は100k(作図時は1M) コンデンサの単位は100n(作図時は1μ)

.include 'LMC6482A.LIB'

.global vcc vee
vcc vcc 0 5
vee vee 0 -5

.ic v(1)=0v
.ic v(4)=3v
.ic v(7)=0v

x1 10 109 intAmp
x2 3 111 intAmp
x3 6 113 intAmp
x4 1 110 invAmp
x5 4 112 invAmp

v1 8 0 1
v2 0 9 2

r1 1 102 100k ;1/Σu
r2 5 103 100k
r3 7 104 100k
r4 7 105 100k ;1/Σp
r5 8 107 33k ;1/vp
* r5 8 107 100k ;1/vp
r6 9 108 100k
r7 2 101 r='50000 / v(4)' ;1/g'
r8 8 106 r='100000 / v(4) / v(4)' ;1/g

* 消費電力プロット用のダミー電圧源
vd1 101 3 0
vd2 102 10 0
vd3 103 6 0
vd4 104 3 0
vd5 105 6 0
vd6 106 10 0
vd7 107 6 0
vd8 108 10 0

vd9 109 1 0 ; x1(積分器)の消費電力プロット用のダミー電圧源
vd10 110 2 0 ; x4(反転増幅器)の消費電力プロット用のダミー電圧源
vd11 111 4 0 ; x2(積分器)の消費電力プロット用のダミー電圧源
vd12 112 5 0 ; x5(反転増幅器)の消費電力プロット用のダミー電圧源
vd13 113 7 0 ; x3(積分器)の消費電力プロット用のダミー電圧源


* 積分器
.subckt intAmp in out
.ic v(1)=0v v(out)=0v
r1 in 1 100k
c1 1 out 100n
x1 0 1 vcc vee out LMC6482A/NS ; IN+ IN- VCC VEE OUT
.ends intAmp

* 反転増幅器
.subckt invAmp in out
.ic v(1)=0v v(out)=0v
r1 in 1 100k
r2 1 out 100k
x1 0 1 vcc vee out LMC6482A/NS
.ends invAmp

.tran 100u 2000m
.control
run
plot v(4) ;φ
plot i(vd1)*(v(2)-v(3)) + i(vd2)*(v(1)-v(10)) + i(vd3)*(v(5)-v(6)) + i(vd4)*(v(7)-v(3)) + i(vd5)*(v(7)-v(6)) + i(vd6)*(v(8)-v(10)) + i(vd7)*(v(8)-v(6)) + i(vd8)*(v(9)-v(10))
+    + i(vd9)*(v(109)-v(10)) + i(vd10)*(v(110)-v(1)) + i(vd11)*(v(111)-v(3)) + i(vd12)*(v(112)-v(4)) + i(vd13)*(v(113)-v(6))
.endc



.end

* DEMO CIRCUIT
* * 関数g(φ)がφ^2 抵抗の単位は100k(作図時は1M) コンデンサの単位は100n(作図時は1μ)

* .include 'LMC6482A.LIB'

* .global vcc vee
* vcc vcc 0 5
* vee vee 0 -5

* .ic v(1)=0v
* .ic v(4)=3v
* .ic v(7)=0v

* x1 10 1 intAmp
* x2 3 4 intAmp
* x3 6 7 intAmp
* x4 1 2 invAmp
* x5 4 5 invAmp

* v1 8 0 1
* v2 0 9 2

* r1 1 10 100k ;1/Σu
* r2 5 6 100k
* r3 7 3 100k
* r4 7 6 100k ;1/Σp
* r5 8 6 33k ;1/vp
* r6 9 10 100k
* r7 2 3 r='50000 / v(4)' ;1/g'
* r8 8 10 r='100000 / v(4) / v(4)' ;1/g

* * 積分器
* .subckt intAmp in out
* .ic v(1)=0v v(out)=0v
* r1 in 1 100k
* c1 1 out 100n
* x1 0 1 vcc vee out LMC6482A/NS ; IN+ IN- VCC VEE OUT
* .ends intAmp

* * 反転増幅器
* .subckt invAmp in out
* .ic v(1)=0v v(out)=0v
* r1 in 1 100k
* r2 1 out 100k
* x1 0 1 vcc vee out LMC6482A/NS
* .ends invAmp

* .tran 100u 2000m
* .control
* run
* plot v(4) ;φ
* .endc

* .end

